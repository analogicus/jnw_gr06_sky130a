magic
tech sky130A
magscale 1 2
timestamp 1742994806
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0
timestamp 1742994806
transform 1 0 1152 0 1 4800
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1742994806
transform 1 0 1152 0 1 4000
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1742994806
transform 1 0 1152 0 1 3198
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1742994806
transform 1 0 1152 0 1 1600
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1742994806
transform 1 0 1152 0 1 800
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1742994806
transform 1 0 1152 0 1 0
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  xa2
timestamp 1742994806
transform 1 0 -762 0 1 0
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  xa3
timestamp 1742994806
transform 1 0 -760 0 1 800
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  xb5[3:0]
timestamp 1742994806
transform 1 0 1152 0 1 2400
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  xb6[3:0]
timestamp 1742994806
transform 1 0 1152 0 1 5600
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  xc6
timestamp 1742994806
transform 1 0 4800 0 1 -8
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  xc7
timestamp 1742994806
transform 1 0 4798 0 1 800
box 0 -1200 361 200
use JNWTR_RPPO16  xd5 ../JNW_TR_SKY130A
timestamp 1742987017
transform 1 0 3420 0 1 2446
box 0 0 4472 3440
use JNWTR_RPPO16  xe4
timestamp 1742987017
transform 1 0 8070 0 1 410
box 0 0 4472 3440
use JNWTR_RPPO16  xf3
timestamp 1742987017
transform 1 0 12870 0 1 1376
box 0 0 4472 3440
<< properties >>
string FIXED_BBOX 0 0 16872 3440
<< end >>
