magic
tech sky130A
magscale 1 2
timestamp 1743333401
<< locali >>
rect 13954 16234 14146 16500
rect 17364 16590 21646 16702
rect 15106 16234 15298 16500
rect 22730 16438 22970 16698
rect 17682 16166 17818 16406
rect 18468 16166 18608 16406
rect 19812 16182 19954 16422
rect 20624 16182 20764 16422
rect 21936 16198 22070 16438
rect 22730 16198 22888 16438
rect 23442 13224 23682 13230
rect 23442 12996 23448 13224
rect 23676 12996 23682 13224
rect 23442 11830 23682 12996
rect 17634 11590 23682 11830
rect 15826 8824 16018 9184
rect 16978 8824 17170 9178
rect 10028 7860 10220 8226
rect 11360 8226 11372 8418
rect 11180 7860 11372 8226
rect 11728 6882 11920 7226
rect 12880 6882 13072 7226
rect 11728 6876 13426 6882
rect 11728 6702 12118 6876
rect 11736 6696 12118 6702
rect 12298 6696 13426 6876
rect 11736 6690 13426 6696
rect 13234 6336 13426 6690
rect 13942 6364 14134 7224
rect 14326 6996 14518 7002
rect 14326 6816 14332 6996
rect 14512 6816 14518 6996
rect 14326 6346 14518 6816
rect 15094 6304 15286 7224
rect 17634 6332 17874 11590
rect 13710 5944 13856 6184
rect 14528 5944 14668 6184
rect 15654 5942 15800 6182
rect 17326 5928 17460 6168
rect 12310 5396 12502 5406
rect 11546 5204 12502 5396
rect 11158 4738 11350 4978
rect 12310 4738 12502 5204
rect 14996 3132 15108 3152
rect 14996 3020 15310 3132
rect 14732 2822 14895 2880
rect 14996 2822 15108 3020
rect 13262 2800 13420 2804
rect 8808 1512 9034 1538
rect 9860 1512 10086 1532
rect 8808 1334 10086 1512
rect 8808 491 9034 1334
rect 9860 491 10086 1334
rect 12228 491 12386 2800
rect 4905 438 9037 491
rect 9855 438 12386 491
rect 4905 260 12386 438
rect 4905 256 9037 260
rect 9855 256 12386 260
rect 9860 254 10086 256
rect 12228 248 12386 256
rect 13262 2788 13568 2800
rect 13262 252 13692 2788
rect 14584 328 14742 2814
rect 14882 2800 15108 2822
rect 14882 328 15040 2800
rect 14584 270 15040 328
rect 15936 2796 16094 2838
rect 16230 2796 16388 2850
rect 15936 298 16388 2796
rect 15936 286 16252 298
rect 14584 262 14940 270
rect 13410 248 13692 252
rect 13436 236 13692 248
rect 13436 208 13594 236
rect 14678 212 14940 262
rect 16094 244 16252 286
rect 18238 -228 18430 942
rect 18646 636 18814 642
rect 18646 480 18652 636
rect 18808 480 18814 636
rect 18646 -254 18814 480
rect 19262 -294 19454 942
rect 19726 -240 19990 92
<< viali >>
rect 13954 16500 14146 16680
rect 15106 16500 15298 16680
rect 17454 16166 17682 16406
rect 18608 16166 18836 16406
rect 19584 16182 19812 16422
rect 20764 16182 20992 16422
rect 21708 16198 21936 16438
rect 22888 16198 23116 16438
rect 23448 12996 23676 13224
rect 6982 10722 7182 10934
rect 15826 9184 16018 9364
rect 16978 9178 17170 9358
rect 10028 8226 10220 8406
rect 11180 8226 11360 8418
rect 12118 6696 12298 6876
rect 14332 6816 14512 6996
rect 13482 5944 13710 6184
rect 14668 5944 14896 6184
rect 15426 5942 15654 6182
rect 17460 5928 17688 6168
rect 11158 4978 11350 5158
rect 18652 480 18808 636
rect 19726 92 19990 344
<< metal1 >>
rect 13954 17112 14146 17114
rect 8958 17106 15328 17112
rect 8958 16914 16018 17106
rect 8958 16900 15328 16914
rect 6976 10934 7188 10946
rect 8958 10934 9170 16900
rect 13954 16686 14146 16900
rect 13942 16680 14158 16686
rect 13942 16500 13954 16680
rect 14146 16500 14158 16680
rect 13942 16494 14158 16500
rect 14338 16082 14530 16900
rect 15106 16686 15298 16900
rect 15094 16680 15310 16686
rect 15094 16500 15106 16680
rect 15298 16500 15310 16680
rect 15094 16494 15310 16500
rect 15826 16406 16018 16914
rect 21702 16438 21942 16450
rect 20912 16434 21708 16438
rect 19578 16422 19818 16434
rect 17448 16406 17688 16418
rect 15822 16166 17454 16406
rect 17682 16166 17688 16406
rect 6976 10722 6982 10934
rect 7182 10722 9186 10934
rect 6976 10710 7188 10722
rect 8430 8418 8622 10722
rect 10412 8418 10604 8432
rect 11174 8418 11366 8430
rect 8423 8406 11180 8418
rect 8423 8226 10028 8406
rect 10220 8226 11180 8406
rect 11360 8226 11366 8418
rect 8423 8220 10934 8226
rect 6647 6103 6653 6169
rect 6719 6103 6725 6169
rect 4647 5960 4713 5966
rect 6653 5902 6719 6103
rect 4647 5888 4713 5894
rect 8430 5404 8622 8220
rect 10412 7706 10604 8220
rect 11174 8214 11366 8226
rect 10284 7008 10348 7318
rect 10284 6938 10348 6944
rect 10796 6642 10988 7500
rect 11978 7214 12042 15126
rect 11978 7206 12048 7214
rect 11984 6642 12048 7206
rect 12112 6882 12304 15146
rect 12496 7606 12688 14982
rect 14212 8810 14276 15982
rect 14338 8486 14530 15890
rect 14212 8052 14276 8292
rect 14724 8092 14916 16156
rect 15826 9626 16018 16166
rect 17448 16154 17688 16166
rect 18602 16406 18842 16418
rect 18982 16406 19584 16422
rect 18602 16166 18608 16406
rect 18836 16182 19584 16406
rect 19812 16182 19818 16422
rect 18836 16166 19374 16182
rect 19578 16170 19818 16182
rect 20758 16422 21708 16434
rect 20758 16182 20764 16422
rect 20992 16198 21708 16422
rect 21936 16198 21942 16438
rect 20992 16182 21570 16198
rect 21702 16186 21942 16198
rect 22882 16438 23122 16450
rect 22882 16198 22888 16438
rect 23116 16198 23682 16438
rect 22882 16186 23122 16198
rect 20758 16170 20998 16182
rect 18602 16154 18842 16166
rect 23442 13230 23682 16198
rect 23436 13224 23688 13230
rect 23436 12996 23448 13224
rect 23676 12996 23688 13224
rect 23436 12990 23688 12996
rect 15820 9434 17170 9626
rect 15826 9370 16018 9434
rect 15814 9364 16030 9370
rect 15814 9184 15826 9364
rect 16018 9184 16030 9364
rect 15814 9178 16030 9184
rect 16210 8672 16402 9434
rect 16978 9364 17170 9434
rect 16966 9358 17182 9364
rect 16966 9178 16978 9358
rect 17170 9178 17182 9358
rect 16966 9172 17182 9178
rect 16082 8092 16146 8330
rect 14724 8052 16146 8092
rect 14212 7988 16146 8052
rect 14724 7900 16146 7988
rect 14724 7430 14916 7900
rect 12106 6876 12310 6882
rect 12106 6696 12118 6876
rect 12298 6696 12310 6876
rect 12106 6690 12310 6696
rect 12496 6664 12688 7346
rect 14198 6664 14262 7212
rect 14326 6996 14518 7380
rect 16594 7284 16786 8504
rect 14326 6816 14332 6996
rect 14512 6816 14518 6996
rect 17352 6892 18558 6956
rect 14326 6804 14518 6816
rect 12496 6642 14286 6664
rect 10796 6472 14286 6642
rect 10796 6456 12688 6472
rect 10804 6450 12688 6456
rect 13476 6184 13716 6196
rect 11930 6051 13482 6184
rect 11698 5985 11704 6051
rect 11770 5985 13482 6051
rect 11926 5944 13482 5985
rect 13710 5944 13716 6184
rect 11158 5404 11350 5406
rect 8430 5212 11736 5404
rect 9612 5114 9804 5212
rect 11158 5164 11350 5212
rect 11542 5204 11736 5212
rect 11146 5158 11362 5164
rect 11146 4978 11158 5158
rect 11350 4978 11362 5158
rect 11146 4972 11362 4978
rect 9612 4916 9804 4922
rect 11542 4580 11734 5204
rect 11926 4640 12118 5944
rect 13476 5932 13716 5944
rect 14662 6184 14902 6196
rect 14662 5944 14668 6184
rect 14896 6182 15230 6184
rect 15420 6182 15660 6194
rect 14896 5944 15426 6182
rect 14662 5942 15426 5944
rect 15654 5942 15660 6182
rect 14662 5932 14902 5942
rect 15420 5930 15660 5942
rect 17454 6168 17694 6180
rect 17454 5928 17460 6168
rect 17688 5928 17694 6168
rect 12015 4607 12081 4640
rect 10496 3244 10560 4052
rect 11416 3848 11480 4222
rect 11544 3762 11736 4480
rect 11416 3244 11480 3382
rect 10496 3180 11480 3244
rect 11416 2944 11480 3180
rect 11416 2874 11480 2880
rect 11928 3119 12120 3614
rect 11928 3053 11999 3119
rect 12065 3053 12120 3119
rect 11928 1168 12120 3053
rect 16600 2550 16840 2552
rect 9612 976 12120 1168
rect 11928 910 12120 976
rect 12464 2548 17196 2550
rect 17454 2548 17694 5928
rect 12464 520 17694 2548
rect 18494 1486 18558 6892
rect 18878 2072 19070 2078
rect 18878 1320 19070 1880
rect 16796 504 17694 520
rect 17454 500 17694 504
rect 18646 636 18814 998
rect 18646 480 18652 636
rect 18808 480 18814 636
rect 18646 468 18814 480
rect 19726 756 19990 762
rect 19726 350 19990 492
rect 19714 344 20002 350
rect 19714 92 19726 344
rect 19990 92 20002 344
rect 19714 86 20002 92
<< via1 >>
rect 6653 6103 6719 6169
rect 4647 5894 4713 5960
rect 10284 6944 10348 7008
rect 11704 5985 11770 6051
rect 9612 4922 9804 5114
rect 11416 2880 11480 2944
rect 11999 3053 12065 3119
rect 18878 1880 19070 2072
rect 19726 492 19990 756
<< metal2 >>
rect 10848 7008 10912 7009
rect 10278 6944 10284 7008
rect 10348 7000 10912 7008
rect 10348 6944 10848 7000
rect 10848 6935 10912 6944
rect 4647 6593 11770 6659
rect 4647 5960 4713 6593
rect 6653 6405 10849 6471
rect 6653 6169 6719 6405
rect 6653 6097 6719 6103
rect 4641 5894 4647 5960
rect 4713 5894 4719 5960
rect 9606 4922 9612 5114
rect 9804 4922 9810 5114
rect 9612 4782 9804 4922
rect 9612 4591 9804 4600
rect 10783 3119 10849 6405
rect 11704 6051 11770 6593
rect 11704 5979 11770 5985
rect 10783 3053 11999 3119
rect 12065 3053 12071 3119
rect 11103 2880 11112 2944
rect 11168 2880 11416 2944
rect 11480 2880 11486 2944
rect 18878 2480 19070 2489
rect 18878 2072 19070 2298
rect 18872 1880 18878 2072
rect 19070 1880 19076 2072
rect 19726 1144 19990 1153
rect 19726 756 19990 890
rect 19720 492 19726 756
rect 19990 492 19996 756
<< via2 >>
rect 10848 6944 10912 7000
rect 9612 4600 9804 4782
rect 11112 2880 11168 2944
rect 18878 2298 19070 2480
rect 19726 890 19990 1144
<< metal3 >>
rect 10843 7000 10917 7005
rect 10843 6944 10848 7000
rect 10912 6944 10917 7000
rect 10843 6939 10917 6944
rect 9607 4782 9809 4787
rect 9607 4600 9612 4782
rect 9804 4600 9809 4782
rect 9607 4595 9809 4600
rect 9612 3536 9804 4595
rect 10848 2944 10912 6939
rect 11107 2944 11173 2949
rect 10772 2880 10778 2944
rect 10842 2880 11112 2944
rect 11168 2880 11173 2944
rect 10848 2874 10912 2880
rect 11107 2875 11173 2880
rect 18878 2485 19070 3876
rect 18873 2480 19075 2485
rect 18873 2298 18878 2480
rect 19070 2298 19075 2480
rect 18873 2293 19075 2298
rect 19726 1604 19990 1610
rect 19726 1149 19990 1342
rect 19721 1144 19995 1149
rect 19721 890 19726 1144
rect 19990 890 19995 1144
rect 19721 885 19995 890
<< via3 >>
rect 10778 2880 10842 2944
rect 19726 1342 19990 1604
<< metal4 >>
rect 10777 2944 10843 2945
rect 10042 2880 10778 2944
rect 10842 2880 10843 2944
rect 10777 2879 10843 2880
rect 19726 1605 19990 4816
rect 19725 1604 19991 1605
rect 19725 1342 19726 1604
rect 19990 1342 19991 1604
rect 19725 1341 19991 1342
use JNWATR_NCH_2C1F2  JNWATR_NCH_2C1F2_0 JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 18334 0 1 790
box -184 -128 1208 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 11826 0 1 9524
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1734044400
transform 1 0 11816 0 1 13576
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1734044400
transform 1 0 11822 0 1 11152
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1734044400
transform 1 0 11820 0 1 10326
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1734044400
transform 1 0 11824 0 1 8698
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_5
timestamp 1734044400
transform 1 0 11826 0 1 7900
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_6
timestamp 1734044400
transform 1 0 14038 0 1 7072
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_7
timestamp 1734044400
transform 1 0 11818 0 1 14402
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_8
timestamp 1734044400
transform 1 0 11822 0 1 12776
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_9
timestamp 1734044400
transform 1 0 11820 0 1 11950
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_10
timestamp 1734044400
transform 1 0 11824 0 1 7074
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 JNW_ATR_SKY130A
timestamp 1743267721
transform 1 0 11256 0 1 3266
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1743267721
transform 1 0 14052 0 1 8176
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1743267721
transform 1 0 11254 0 1 4090
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1743267721
transform 1 0 14048 0 1 9008
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1743267721
transform 1 0 15922 0 1 8176
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1743267721
transform 1 0 14046 0 1 13124
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_6
timestamp 1743267721
transform 1 0 14054 0 1 13956
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_7
timestamp 1743267721
transform 1 0 14052 0 1 9834
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_8
timestamp 1743267721
transform 1 0 14050 0 1 10666
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_9
timestamp 1743267721
transform 1 0 14046 0 1 11492
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_10
timestamp 1743267721
transform 1 0 14050 0 1 12324
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_11
timestamp 1743267721
transform 1 0 14046 0 1 14754
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_12
timestamp 1743267721
transform 1 0 14050 0 1 15586
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_13
timestamp 1743267721
transform 1 0 10124 0 1 7212
box -184 -128 1336 928
use JNWTR_CAPX1  JNWTR_CAPX1_0 JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 9230 0 1 2624
box 0 0 1080 1080
use JNWTR_RPPO4  JNWTR_RPPO4_0 JNW_TR_SKY130A
timestamp 1743265964
transform 1 0 13252 0 1 3024
box 0 0 1880 3440
use JNWTR_RPPO8  JNWTR_RPPO8_0 JNW_TR_SKY130A
timestamp 1743265964
transform 1 0 15206 0 1 3008
box 0 0 2744 3440
use OTA  OTA_0
timestamp 1743272310
transform 1 0 0 0 1 480
box 0 -480 10506 10458
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1734020192
transform 1 0 14832 0 1 1564
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1734020192
transform 1 0 8776 0 1 230
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1734020192
transform 1 0 12132 0 1 186
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1734020192
transform 1 0 13480 0 1 186
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1734020192
transform 1 0 14830 0 1 186
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1734020192
transform 1 0 16178 0 1 186
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1734020192
transform 1 0 12132 0 1 1566
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1734020192
transform 1 0 13476 0 1 1566
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1734020192
transform 1 0 16180 0 1 1562
box 0 0 1340 1340
<< labels >>
flabel space 4890 256 9062 491 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 7182 10722 9186 10934 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal1 16594 7284 16786 7476 0 FreeSans 1600 0 0 0 OUT
port 13 nsew
<< end >>
