magic
tech sky130A
magscale 1 2
timestamp 1743293941
<< locali >>
rect 9694 25080 10082 25192
rect 10174 24916 10558 24928
rect 10414 24688 10558 24916
rect 11230 24688 11380 24928
rect 9970 21570 10082 21896
rect 10378 21190 10526 21430
rect 11192 21190 11340 21430
rect 9938 18068 10050 18398
rect 9916 17694 10502 17934
rect 11174 17694 11308 17934
rect 9964 14806 10076 14902
rect 9964 14624 10076 14680
rect 10374 14384 11996 14690
rect 11044 10664 11236 10974
rect 12068 10784 12260 11022
rect 12068 10664 12700 10784
rect 11044 10644 12700 10664
rect 11044 10488 11434 10644
rect 11590 10592 12700 10644
rect 11590 10488 12461 10592
rect 450 8220 685 8763
rect 11044 8663 12461 10488
rect 8827 8461 12461 8663
rect 11044 8220 12461 8461
rect 450 7985 12511 8220
rect 11044 7188 12461 7985
<< viali >>
rect 17764 25252 17964 25464
rect 9594 25080 9694 25192
rect 10174 24688 10414 24916
rect 11380 24688 11608 24928
rect 10150 21190 10378 21430
rect 11340 21190 11568 21430
rect 11308 17694 11536 17934
rect 11434 10488 11590 10644
rect 12700 10592 12880 10784
<< metal1 >>
rect 1544 25560 1756 25800
rect 10671 25560 11045 26821
rect 1544 25476 17918 25560
rect 1544 25464 17970 25476
rect 1544 25348 17764 25464
rect 1544 25172 1756 25348
rect 7275 25252 17764 25348
rect 17964 25252 17970 25464
rect 7275 25192 11618 25252
rect 17758 25240 17970 25252
rect 7275 25186 9594 25192
rect 8438 25080 9594 25186
rect 9694 25186 11618 25192
rect 9694 25080 9700 25186
rect 9588 25068 9700 25080
rect 11374 24928 11614 25186
rect 10162 24916 10426 24922
rect 10162 24688 10174 24916
rect 10414 24688 10426 24916
rect 10162 24682 10426 24688
rect 11374 24688 11380 24928
rect 11608 24688 11614 24928
rect 10174 21868 10414 24682
rect 11374 24676 11614 24688
rect 10174 21628 11574 21868
rect 10144 21430 10384 21442
rect 10144 21190 10150 21430
rect 10378 21190 10384 21430
rect 10144 19729 10384 21190
rect 11334 21430 11574 21628
rect 11334 21190 11340 21430
rect 11568 21190 11574 21430
rect 11334 21178 11574 21190
rect 18519 20498 18585 20504
rect 10144 19663 10631 19729
rect 10697 19663 10703 19729
rect 10144 18334 10384 19663
rect 16527 19305 16593 20490
rect 18519 20426 18585 20432
rect 16527 19233 16593 19239
rect 22204 18390 22900 18582
rect 10134 18094 11542 18334
rect 11302 17934 11542 18094
rect 11302 17694 11308 17934
rect 11536 17694 11542 17934
rect 11302 17682 11542 17694
rect 9128 15748 9320 15754
rect 9128 15550 9320 15556
rect 10780 11960 11364 12024
rect 11300 11454 11364 11960
rect 11684 11844 11876 11850
rect 11684 11254 11876 11652
rect 12694 11386 12886 11392
rect 11428 10644 11596 11030
rect 11428 10488 11434 10644
rect 11590 10488 11596 10644
rect 12694 10784 12886 11194
rect 12694 10592 12700 10784
rect 12880 10592 12886 10784
rect 12694 10580 12886 10592
rect 11428 10476 11596 10488
<< via1 >>
rect 10631 19663 10697 19729
rect 18519 20432 18585 20498
rect 16527 19239 16593 19305
rect 9128 15556 9320 15748
rect 11684 11652 11876 11844
rect 12694 11194 12886 11386
<< metal2 >>
rect 18513 20432 18519 20498
rect 18585 20432 18591 20498
rect 10631 19729 10697 19735
rect 18519 19729 18585 20432
rect 10697 19663 18585 19729
rect 10631 19657 10697 19663
rect 16521 19239 16527 19305
rect 16593 19239 16599 19305
rect 9122 15556 9128 15748
rect 9320 15556 9326 15748
rect 9128 15523 9320 15556
rect 16527 15523 16593 19239
rect 9128 15457 16593 15523
rect 9128 15234 9320 15457
rect 9128 15043 9320 15052
rect 11684 12242 11876 12251
rect 11684 11844 11876 12060
rect 12694 11990 12886 11999
rect 11678 11652 11684 11844
rect 11876 11652 11882 11844
rect 12694 11386 12886 11808
rect 12688 11194 12694 11386
rect 12886 11194 12892 11386
<< via2 >>
rect 9128 15052 9320 15234
rect 11684 12060 11876 12242
rect 12694 11808 12886 11990
<< metal3 >>
rect 9123 15234 9325 15239
rect 9123 15052 9128 15234
rect 9320 15052 9325 15234
rect 9123 15047 9325 15052
rect 9128 13090 9320 15047
rect 9128 13050 11796 13090
rect 9128 12898 11876 13050
rect 11684 12247 11876 12898
rect 12694 12692 12886 12698
rect 11679 12242 11881 12247
rect 11679 12060 11684 12242
rect 11876 12060 11881 12242
rect 11679 12055 11881 12060
rect 12694 11995 12886 12502
rect 12689 11990 12891 11995
rect 12689 11808 12694 11990
rect 12886 11808 12891 11990
rect 12689 11803 12891 11808
<< via3 >>
rect 12694 12502 12886 12692
<< metal4 >>
rect 11970 12924 12886 13116
rect 12694 12693 12886 12924
rect 12693 12692 12887 12693
rect 12693 12502 12694 12692
rect 12886 12502 12887 12692
rect 12693 12501 12887 12502
use JNWATR_PCH_2C1F2  JNWATR_PCH_2C1F2_0 JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 11140 0 1 10822
box -184 -128 1208 928
use JNWTR_CAPX1  JNWTR_CAPX1_0 JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 11172 0 1 12498
box 0 0 1080 1080
use JNWTR_RPPO4  JNWTR_RPPO4_0 JNW_TR_SKY130A
timestamp 1743265964
transform 1 0 9898 0 1 14774
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_1
timestamp 1743265964
transform 1 0 9954 0 1 21768
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_2
timestamp 1743265964
transform 1 0 9922 0 1 18270
box 0 0 1880 3440
use OTA  OTA_1
timestamp 1743272310
transform 1 0 11890 0 1 15010
box 0 -480 10506 10458
use temp_affected_current  temp_affected_current_1
timestamp 1743290148
transform 1 0 -7466 0 1 8272
box 0 0 17950 17114
<< labels >>
flabel metal1 1544 25588 1756 25800 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel locali 450 7985 685 8220 0 FreeSans 1600 0 0 0 VSS
port 13 nsew
flabel metal1 10780 11960 10844 12024 0 FreeSans 1600 0 0 0 reset
port 17 nsew
flabel metal1 22708 18390 22900 18582 0 FreeSans 1600 0 0 0 OUT
port 19 nsew
flabel metal1 10671 26433 11045 26807 0 FreeSans 1600 0 0 0 VDD
port 21 nsew
<< end >>
