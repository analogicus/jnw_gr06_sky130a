magic
tech sky130A
magscale 1 2
timestamp 1743283403
<< locali >>
rect 16406 106 21105 1872
<< metal1 >>
rect 16176 18092 18604 18284
rect 16158 15976 18318 16168
rect 8380 3862 8386 4054
rect 8578 3862 8584 4054
<< via1 >>
rect 8386 3862 8578 4054
<< metal2 >>
rect 8386 4054 8578 4060
rect 8578 3862 8587 4054
rect 8386 3856 8578 3862
<< via2 >>
rect 8396 3862 8578 4054
<< metal3 >>
rect 8387 3857 8393 4059
rect 8583 3857 8589 4059
<< via3 >>
rect 8393 4054 8583 4059
rect 8393 3862 8396 4054
rect 8396 3862 8578 4054
rect 8578 3862 8583 4054
rect 8393 3857 8583 3862
<< metal4 >>
rect 8392 4059 8584 4060
rect 8392 3857 8393 4059
rect 8583 4054 8584 4059
rect 10424 4054 10616 4182
rect 10664 4054 10856 4194
rect 8583 3862 10856 4054
rect 8583 3857 8584 3862
rect 8392 3856 8584 3857
use temp_affected_current  temp_affected_current_1
timestamp 1743272310
transform 1 0 9438 0 1 4970
box -9440 -4968 8788 13334
<< labels >>
flabel locali 19339 106 21105 1872 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal1 18412 18092 18604 18284 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel metal1 18126 15976 18318 16168 0 FreeSans 1600 0 0 0 TEST
port 4 nsew
<< end >>
