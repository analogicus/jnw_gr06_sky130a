    
    *TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/temp_affected_current_lpe.spi
#else
.include ../../../work/xsch/temp_affected_current.spice
#endif


Rout OUT VSS 1k ac=10k m=1

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3 

.temp 27
*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS  dc {AVDD}



*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------


*----------------------------------------------------------------
* SAVES
*----------------------------------------------------------------
.save v(OUT) v(GATE)
.option savecurrents
*.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit


optran 0 0 0 1n 1u 0
dc temp -60 120 1




write
quit


.endc

.end
