magic
tech sky130A
magscale 1 2
timestamp 1743679690
<< locali >>
rect 6258 10454 6450 10458
rect 5874 10434 7224 10454
rect 5872 10262 7224 10434
rect 5872 10242 7218 10262
rect 5874 9404 6066 10242
rect 6258 9848 6450 10242
rect 6258 9668 6264 9848
rect 6444 9668 6450 9848
rect 6258 9662 6450 9668
rect 7026 9358 7218 10242
rect 5878 8284 6070 8852
rect 7030 8288 7222 8908
rect 48 6804 160 7140
rect 4922 7028 5114 7334
rect 6074 7028 6266 7320
rect 6904 7036 7096 7320
rect 8236 7322 8248 7514
rect 8056 7018 8248 7322
rect 28 3300 140 3622
rect 4922 1788 5114 2498
rect 5306 2158 5498 2164
rect 5306 1978 5312 2158
rect 5492 1978 5498 2158
rect 5306 1788 5498 1978
rect 6074 1788 6266 2504
rect 6906 1788 7098 2496
rect 7290 2182 7482 2188
rect 7290 2002 7296 2182
rect 7476 2002 7482 2182
rect 7290 1788 7482 2002
rect 8058 1788 8250 2522
rect 4922 1786 8250 1788
rect 4890 1596 8250 1786
rect 16 -350 128 128
rect 16 -462 28 -350
rect 4890 -246 5130 1596
rect 8058 1592 8250 1596
rect 4890 -474 4896 -246
rect 5124 -474 5130 -246
rect 4890 -480 5130 -474
<< viali >>
rect 396 9932 636 10160
rect 3912 9932 4140 10172
rect 6264 9668 6444 9848
rect 4922 7334 5114 7514
rect 6074 7320 6266 7500
rect 6904 7320 7096 7500
rect 8056 7322 8236 7514
rect 376 6414 604 6654
rect 3874 6420 4102 6648
rect 364 2920 604 3148
rect 3866 2928 4094 3156
rect 5312 1978 5492 2158
rect 7296 2002 7476 2182
rect 28 -462 128 -350
rect 4896 -474 5124 -246
<< metal1 >>
rect 3906 10172 4146 10184
rect 6642 10172 6834 10174
rect 384 10160 648 10166
rect 384 9932 396 10160
rect 636 9932 648 10160
rect 384 9926 648 9932
rect 3906 9932 3912 10172
rect 4140 9932 6834 10172
rect 396 7638 636 9926
rect 3906 9920 4146 9932
rect 6130 9406 6194 9932
rect 6258 9848 6450 9860
rect 6258 9668 6264 9848
rect 6444 9668 6450 9848
rect 6258 9220 6450 9668
rect 6642 9292 6834 9932
rect 6134 8304 6198 8928
rect 6262 8128 6454 9018
rect 396 7398 4108 7638
rect 370 6654 610 6666
rect 370 6414 376 6654
rect 604 6414 610 6654
rect 370 5198 610 6414
rect 3868 6648 4108 7398
rect 4910 7514 5612 7520
rect 4910 7334 4922 7514
rect 5114 7510 5612 7514
rect 6646 7510 6838 7922
rect 8050 7514 8242 7526
rect 7146 7510 8056 7514
rect 5114 7500 8056 7510
rect 5114 7334 6074 7500
rect 4910 7328 6074 7334
rect 5306 7320 6074 7328
rect 6266 7320 6904 7500
rect 7096 7322 8056 7500
rect 8236 7322 8242 7514
rect 7096 7320 7486 7322
rect 5306 7318 7486 7320
rect 5306 6780 5498 7318
rect 6062 7314 6278 7318
rect 6892 7314 7108 7318
rect 7294 6880 7486 7318
rect 8050 7310 8242 7322
rect 3868 6420 3874 6648
rect 4102 6420 4108 6648
rect 3868 6408 4108 6420
rect 5178 5480 5242 6486
rect 4637 5414 5242 5480
rect 370 4958 4100 5198
rect 3860 3156 4100 4958
rect 5178 4538 5242 5414
rect 5306 4284 5498 6684
rect 5688 4384 5880 6686
rect 7160 5488 7224 6500
rect 6619 5422 7224 5488
rect 7160 4572 7224 5422
rect 7286 4328 7478 6640
rect 7672 4360 7864 6716
rect 5688 3502 5880 4172
rect 7670 3572 7862 4178
rect 352 3148 616 3154
rect 352 2920 364 3148
rect 604 2920 616 3148
rect 352 2914 616 2920
rect 3860 2928 3866 3156
rect 4094 2928 4100 3156
rect 5178 3492 5896 3502
rect 5178 3438 7226 3492
rect 5178 3020 5242 3438
rect 5688 3428 7226 3438
rect 3860 2916 4100 2928
rect 364 -240 604 2914
rect 5688 2706 5880 3428
rect 7162 2964 7226 3428
rect 7670 3380 10506 3572
rect 7670 2730 7862 3380
rect 5306 2158 5498 2650
rect 5306 1978 5312 2158
rect 5492 1978 5498 2158
rect 7290 2182 7482 2648
rect 7290 2002 7296 2182
rect 7476 2002 7482 2182
rect 7290 1990 7482 2002
rect 5306 1966 5498 1978
rect 364 -246 5136 -240
rect 22 -350 134 -338
rect 364 -350 4896 -246
rect 22 -462 28 -350
rect 128 -462 4896 -350
rect 22 -474 134 -462
rect 364 -474 4896 -462
rect 5124 -474 5136 -246
rect 364 -480 5136 -474
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 5018 0 1 2346
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1734044400
transform 1 0 7002 0 1 2344
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 JNW_ATR_SKY130A
timestamp 1743267721
transform 1 0 6998 0 1 4728
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1743267721
transform 1 0 6998 0 1 3906
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1743267721
transform 1 0 7000 0 1 5566
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1743267721
transform 1 0 7000 0 1 6388
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1743267721
transform 1 0 5016 0 1 3898
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1743267721
transform 1 0 5016 0 1 4720
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_6
timestamp 1743267721
transform 1 0 5018 0 1 5558
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_7
timestamp 1743267721
transform 1 0 5018 0 1 6380
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_8
timestamp 1743267721
transform 1 0 5972 0 1 7790
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_9
timestamp 1743267721
transform 1 0 5968 0 1 8794
box -184 -128 1336 928
use JNWTR_RPPO16  JNWTR_RPPO16_0 JNW_TR_SKY130A
timestamp 1743679690
transform 1 0 12 0 1 3494
box 0 0 4472 3440
use JNWTR_RPPO16  JNWTR_RPPO16_1
timestamp 1743679690
transform 1 0 0 0 1 0
box 0 0 4472 3440
use JNWTR_RPPO16  JNWTR_RPPO16_3
timestamp 1743679690
transform 1 0 32 0 1 7012
box 0 0 4472 3440
<< labels >>
flabel metal1 364 -480 604 2920 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 4637 5414 5242 5480 0 FreeSans 1600 0 0 0 IN+
port 9 nsew
flabel metal1 6619 5422 7224 5488 0 FreeSans 1600 0 0 0 IN-
port 11 nsew
flabel locali 5874 10242 7218 10454 0 FreeSans 1600 0 0 0 VDD
port 13 nsew
flabel metal1 7670 3380 10506 3572 0 FreeSans 1600 0 0 0 OUT
port 15 nsew
<< end >>
