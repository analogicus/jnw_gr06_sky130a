magic
tech sky130A
magscale 1 2
timestamp 1742943600
<< checkpaint >>
rect 0 0 11448 1080
use JNWATR_PCH_4C5F0 x1 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 0
box 0 0 1152 800
use JNWATR_PCH_4C5F0 x2 ../JNW_ATR_SKY130A
transform 1 0 1152 0 1 0
box 1152 0 2304 800
use OTA x3 ../JNW_GR06_SKY130A
transform 1 0 2304 0 1 0
box 2304 0 4608 800
use JNWATR_PCH_4C5F0 x4 ../JNW_ATR_SKY130A
transform 1 0 4608 0 1 0
box 4608 0 5760 800
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 0
box 5760 0 6912 800
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 800
box 5760 800 6912 1600
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 1600
box 5760 1600 6912 2400
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 2400
box 5760 2400 6912 3200
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 3200
box 5760 3200 6912 4000
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 4000
box 5760 4000 6912 4800
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 4800
box 5760 4800 6912 5600
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 5600
box 5760 5600 6912 6400
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 6400
box 5760 6400 6912 7200
use JNWATR_NCH_4C5F0 x5[9:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 7200
box 5760 7200 6912 8000
use JNWATR_NCH_4C5F0 x6 ../JNW_ATR_SKY130A
transform 1 0 6912 0 1 0
box 6912 0 8064 800
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 0
box 8064 0 9216 800
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 800
box 8064 800 9216 1600
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 1600
box 8064 1600 9216 2400
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 2400
box 8064 2400 9216 3200
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 3200
box 8064 3200 9216 4000
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 4000
box 8064 4000 9216 4800
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 4800
box 8064 4800 9216 5600
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 5600
box 8064 5600 9216 6400
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 6400
box 8064 6400 9216 7200
use JNWATR_PCH_4C5F0 x7[9:0] ../JNW_ATR_SKY130A
transform 1 0 8064 0 1 7200
box 8064 7200 9216 8000
use JNWTR_CAPX1 x8 ../JNW_TR_SKY130A
transform 1 0 9216 0 1 0
box 9216 0 10296 1080
use JNWATR_PCH_4C5F0 x9 ../JNW_ATR_SKY130A
transform 1 0 10296 0 1 0
box 10296 0 11448 800
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 11448 1080
<< end >>
