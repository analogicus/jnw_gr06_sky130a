magic
tech sky130A
magscale 1 2
timestamp 1743272310
<< locali >>
rect 1446 12824 1638 13122
rect 2778 13122 2790 13314
rect 2598 12824 2790 13122
rect 3686 12798 3878 13130
rect 4838 12798 5030 13134
rect 5952 12776 6144 13136
rect 7284 13130 7296 13322
rect 7104 12776 7296 13130
rect 2620 3786 2632 3794
rect 2696 3786 2812 3794
rect 1468 3418 1660 3784
rect 1844 3420 2586 3426
rect 1844 3418 1850 3420
rect 1468 3232 1850 3418
rect 2038 3418 2586 3420
rect 2620 3418 2812 3786
rect 3674 3418 3866 3750
rect 4058 3418 4596 3422
rect 4826 3418 5018 3750
rect 2038 3416 5018 3418
rect 2038 3236 4064 3416
rect 4244 3236 5018 3416
rect 2038 3232 5018 3236
rect 1468 3230 5018 3232
rect 1476 3226 4998 3230
rect 3674 3218 3866 3226
rect 7372 2376 8162 2616
rect -96 1472 96 1842
rect 1056 1472 1248 1832
rect 7922 -444 8162 2376
rect 3308 -642 8162 -444
rect 8546 -642 8734 -626
rect 3308 -730 8734 -642
rect 3302 -826 8734 -730
rect 3302 -1730 3516 -826
rect 4366 -1730 4908 -826
rect 5764 -1730 6306 -826
rect 7160 -1730 7702 -826
rect 8546 -1730 8734 -826
rect 3302 -1878 8734 -1730
rect 618 -2234 1908 -2000
rect 3302 -2042 8762 -1878
rect 3302 -2226 8766 -2042
rect 646 -3058 848 -2234
rect 1692 -3058 1902 -2234
rect 646 -3212 1902 -3058
rect 3302 -3098 3516 -2226
rect 4366 -3098 4908 -2226
rect 5764 -3098 6306 -2226
rect 7160 -3098 7702 -2226
rect 8546 -3098 8734 -2226
rect 3302 -3212 8746 -3098
rect -4476 -3282 8746 -3212
rect -4476 -4864 8734 -3282
rect -4476 -4870 4300 -4864
<< viali >>
rect 1446 13122 1638 13302
rect 2598 13122 2778 13314
rect 3686 13130 3878 13310
rect 4838 13134 5030 13314
rect 5952 13136 6144 13316
rect 7104 13130 7284 13322
rect -2422 5754 -2222 5966
rect 1850 3232 2038 3420
rect 4064 3236 4244 3416
rect 3654 2366 3882 2606
rect 4578 2366 4806 2606
rect 5548 2372 5776 2600
rect -96 1842 96 2022
rect 1056 1832 1248 2012
<< metal1 >>
rect 2592 13314 2784 13326
rect 7098 13322 7290 13334
rect 3674 13314 3890 13316
rect 4826 13314 5042 13320
rect 5640 13316 6156 13322
rect 5640 13314 5952 13316
rect -119 13308 308 13313
rect 1036 13308 2598 13314
rect -142 13302 2598 13308
rect -142 13122 1446 13302
rect 1638 13122 2598 13302
rect 2778 13310 4838 13314
rect 2778 13130 3686 13310
rect 3878 13134 4838 13310
rect 5030 13136 5952 13314
rect 6144 13314 6156 13316
rect 7098 13314 7104 13322
rect 6144 13136 7104 13314
rect 5030 13134 7104 13136
rect 3878 13130 7104 13134
rect 7284 13314 7290 13322
rect 7284 13130 7296 13314
rect 2778 13122 7296 13130
rect -142 13116 1650 13122
rect -119 6011 308 13116
rect 1830 12672 2022 13122
rect 2592 13110 2784 13122
rect 838 12216 1766 12280
rect 844 11708 908 12216
rect 2228 12002 2428 12544
rect 1716 11930 2428 12002
rect 1716 11740 1788 11930
rect 844 11638 908 11644
rect -2409 5978 318 6011
rect -2428 5966 318 5978
rect -2428 5754 -2422 5966
rect -2222 5754 318 5966
rect -2428 5742 318 5754
rect -2409 5584 318 5742
rect -109 2449 318 5584
rect 1724 4294 1788 11740
rect 1844 3924 2036 11696
rect 2228 11618 2428 11930
rect 2236 4210 2428 11618
rect 3952 5352 4016 12854
rect 3952 4596 4016 4830
rect 4070 4770 4262 13122
rect 4464 12807 4656 12902
rect 4454 12605 6263 12807
rect 6336 12624 6528 13122
rect 7098 13118 7290 13122
rect 4464 4596 4656 12605
rect 6720 10984 6912 12382
rect 3952 4532 4656 4596
rect 2236 4146 3994 4210
rect 1844 3420 2044 3924
rect 2236 3752 2428 4146
rect 1844 3232 1850 3420
rect 2038 3232 2044 3420
rect 1844 3220 2044 3232
rect 4058 3416 4250 3924
rect 4464 3648 4656 4532
rect 4058 3236 4064 3416
rect 4244 3236 4250 3416
rect 4058 3224 4250 3236
rect 3648 2606 3888 2618
rect -109 2440 2196 2449
rect -112 2083 2196 2440
rect 2826 2366 3654 2606
rect 3882 2366 3888 2606
rect -112 2071 1818 2083
rect -112 2028 1246 2071
rect -112 2022 1264 2028
rect -112 1842 -96 2022
rect 96 2012 1264 2022
rect 96 1842 1056 2012
rect -112 1832 1056 1842
rect 1248 1836 1264 2012
rect 1248 1832 1260 1836
rect -112 1828 1260 1832
rect -4840 1392 -4834 1584
rect -4642 1392 -4636 1584
rect -4834 1118 -4642 1392
rect 288 1306 480 1828
rect 1044 1826 1260 1828
rect 1812 1705 1818 2071
rect 2196 1705 2202 2083
rect 672 1584 864 1590
rect 672 1386 864 1392
rect 2826 1166 3090 2366
rect 3648 2354 3888 2366
rect 4572 2606 4812 2618
rect 4572 2366 4578 2606
rect 4806 2600 5788 2606
rect 4806 2372 5548 2600
rect 5776 2372 5788 2600
rect 4806 2366 5788 2372
rect 4572 2354 4812 2366
rect -4834 926 -4202 1118
rect -2814 -432 -2622 1010
rect 160 840 224 946
rect 158 678 224 840
rect 158 120 222 678
rect 288 332 480 1164
rect 672 974 3090 1166
rect 672 270 864 368
rect 158 -216 224 120
rect -2814 -630 -2622 -624
rect -734 -280 224 -216
rect -734 -784 -670 -280
rect 160 -294 224 -280
rect 672 78 1458 270
rect 672 -432 864 78
rect 672 -632 864 -624
rect -560 -784 -496 -778
rect -734 -848 -560 -784
rect -560 -854 -496 -848
rect 1266 -2660 1458 78
<< via1 >>
rect 844 11644 908 11708
rect -4834 1392 -4642 1584
rect 1818 1705 2196 2083
rect 672 1392 864 1584
rect -2814 -624 -2622 -432
rect 672 -624 864 -432
rect -560 -848 -496 -784
<< metal2 >>
rect 838 11644 844 11708
rect 908 11644 914 11708
rect 844 10730 908 11644
rect 844 10665 908 10674
rect 1818 2083 2196 2089
rect 1814 1710 1818 2078
rect 2196 1710 2200 2078
rect 1818 1699 2196 1705
rect -4834 1584 -4642 1590
rect -4642 1392 672 1584
rect 864 1392 870 1584
rect -4834 1386 -4642 1392
rect -2820 -624 -2814 -432
rect -2622 -624 672 -432
rect 864 -624 870 -432
rect -264 -784 -208 -779
rect -566 -848 -560 -784
rect -496 -788 -204 -784
rect -496 -844 -264 -788
rect -208 -844 -204 -788
rect -496 -848 -204 -844
rect -264 -853 -208 -848
<< via2 >>
rect 844 10674 908 10730
rect 1823 1710 2191 2078
rect -264 -844 -208 -788
<< metal3 >>
rect 839 10730 913 10735
rect 839 10674 844 10730
rect 908 10674 913 10730
rect 839 10669 913 10674
rect 844 9790 908 10669
rect 844 9720 908 9726
rect 1818 2078 2196 2083
rect 1818 1710 1823 2078
rect 2191 1710 2196 2078
rect 1818 -394 2196 1710
rect -269 -784 -203 -783
rect -44 -784 20 -778
rect -269 -788 -44 -784
rect -269 -844 -264 -788
rect -208 -844 -44 -788
rect -269 -848 -44 -844
rect -269 -849 -203 -848
rect -44 -854 20 -848
<< via3 >>
rect 844 9726 908 9790
rect -44 -848 20 -784
<< metal4 >>
rect 843 9790 909 9791
rect 843 9726 844 9790
rect 908 9726 909 9790
rect 843 9725 909 9726
rect -45 -784 21 -783
rect 844 -784 908 9725
rect -45 -848 -44 -784
rect 20 -848 1364 -784
rect -45 -849 21 -848
rect 844 -850 908 -848
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 3770 0 1 3598
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1734044400
transform 1 0 1556 0 1 11084
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1734044400
transform 1 0 1562 0 1 5284
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1734044400
transform 1 0 1562 0 1 4462
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1734044400
transform 1 0 1560 0 1 6950
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_5
timestamp 1734044400
transform 1 0 1558 0 1 7788
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_6
timestamp 1734044400
transform 1 0 1558 0 1 10246
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_7
timestamp 1734044400
transform 1 0 1560 0 1 6122
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_8
timestamp 1734044400
transform 1 0 1556 0 1 9448
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_9
timestamp 1734044400
transform 1 0 1558 0 1 8610
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_10
timestamp 1734044400
transform 1 0 1564 0 1 3624
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 JNW_ATR_SKY130A
timestamp 1743267721
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1743267721
transform 1 0 0 0 1 824
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1743267721
transform 1 0 3792 0 1 6372
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1743267721
transform 1 0 1542 0 1 12176
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1743267721
transform 1 0 3790 0 1 7216
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1743267721
transform 1 0 3790 0 1 5570
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_6
timestamp 1743267721
transform 1 0 3792 0 1 4726
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_7
timestamp 1743267721
transform 1 0 3792 0 1 8016
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_8
timestamp 1743267721
transform 1 0 3790 0 1 8860
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_9
timestamp 1743267721
transform 1 0 3786 0 1 11306
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_10
timestamp 1743267721
transform 1 0 3782 0 1 12150
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_11
timestamp 1743267721
transform 1 0 3792 0 1 9662
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_12
timestamp 1743267721
transform 1 0 3790 0 1 10506
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_13
timestamp 1743267721
transform 1 0 6048 0 1 12128
box -184 -128 1336 928
use JNWTR_CAPX1  JNWTR_CAPX1_0 JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 1120 0 1 -1176
box 0 0 1080 1080
use JNWTR_RPPO4  JNWTR_RPPO4_0 JNW_TR_SKY130A
timestamp 1743265964
transform 1 0 3290 0 1 -554
box 0 0 1880 3440
use JNWTR_RPPO8  JNWTR_RPPO8_0 JNW_TR_SKY130A
timestamp 1743265964
transform 1 0 5232 0 1 -544
box 0 0 2744 3440
use OTA  OTA_0
timestamp 1743272310
transform 1 0 -9440 0 1 -4488
box 0 -480 10506 10458
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1734020192
transform 1 0 4664 0 1 -1940
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1734020192
transform 1 0 590 0 1 -3314
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1734020192
transform 1 0 7436 0 1 -1924
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1734020192
transform 1 0 3268 0 1 -1940
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1734020192
transform 1 0 3280 0 1 -3312
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1734020192
transform 1 0 6062 0 1 -1940
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1734020192
transform 1 0 4676 0 1 -3312
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1734020192
transform 1 0 6074 0 1 -3312
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1734020192
transform 1 0 7448 0 1 -3296
box 0 0 1340 1340
<< labels >>
flabel locali -4476 -4870 4300 -3212 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 6720 10984 6912 11176 0 FreeSans 1600 0 0 0 OUT
port 3 nsew
<< end >>
