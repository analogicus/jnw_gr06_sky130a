magic
tech sky130A
magscale 1 2
timestamp 1742994806
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0
timestamp 1742994806
transform 1 0 2232 0 1 7200
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1742994806
transform 1 0 2232 0 1 6400
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1742994806
transform 1 0 2232 0 1 5600
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1742994806
transform 1 0 2232 0 1 4800
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1742994806
transform 1 0 2232 0 1 4000
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_5
timestamp 1742994806
transform 1 0 2232 0 1 3200
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_6
timestamp 1742994806
transform 1 0 2232 0 1 2400
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_7
timestamp 1742994806
transform 1 0 2232 0 1 1600
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_8
timestamp 1742994806
transform 1 0 2232 0 1 800
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0
timestamp 1742994806
transform 1 0 0 0 1 8800
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1742994806
transform 1 0 0 0 1 8000
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1742994806
transform 1 0 0 0 1 7200
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1742994806
transform 1 0 0 0 1 6400
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1742994806
transform 1 0 0 0 1 5600
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1742994806
transform 1 0 0 0 1 4800
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_6
timestamp 1742994806
transform 1 0 0 0 1 4000
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_7
timestamp 1742994806
transform 1 0 0 0 1 3200
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_8
timestamp 1742994806
transform 1 0 0 0 1 2400
box 0 -1200 361 200
use JNWTR_RPPO4  JNWTR_RPPO4_0 JNW_TR_SKY130A
timestamp 1742990092
transform 1 0 4868 0 1 136
box 0 0 1880 3440
use JNWATR_PCH_4C5F0  xa1
timestamp 1742994806
transform 1 0 0 0 1 0
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  xa2
timestamp 1742994806
transform 1 0 0 0 1 800
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  xa4
timestamp 1742994806
transform 1 0 0 0 1 1600
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  xa5[9:0]
timestamp 1742994806
transform 1 0 0 0 1 9600
box 0 -1200 361 200
use JNWATR_PCH_4C5F0  xa9
timestamp 1742994806
transform 1 0 0 0 1 10400
box 0 -1200 361 200
use JNWTR_CAPX1  xb8 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 4720 0 1 3870
box 0 0 1080 1080
use JNWATR_NCH_4C5F0  xc1[9:0]
timestamp 1742994806
transform 1 0 2232 0 1 8000
box 0 -1200 361 200
use JNWATR_NCH_4C5F0  xc11
timestamp 1742994806
transform 1 0 2232 0 1 0
box 0 -1200 361 200
use JNWTR_RPPO8  xd7 ../JNW_TR_SKY130A
timestamp 1742990092
transform 1 0 4748 0 1 5674
box 0 0 2744 3440
use OTA  xe3
timestamp 1742994806
transform 1 0 8602 0 1 -158
box -762 -1208 17342 5886
<< properties >>
string FIXED_BBOX 0 0 23000 11200
<< end >>
