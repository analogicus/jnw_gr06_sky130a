magic
tech sky130A
magscale 1 2
timestamp 1743030000
<< checkpaint >>
rect 0 0 16952 7480
use JNWATR_PCH_4C5F0 x1 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 0
box 0 0 1152 800
use JNWATR_PCH_4C5F0 x2 ../JNW_ATR_SKY130A
transform 1 0 1832 0 1 0
box 1832 0 2984 800
use JNWTR_RPPO16 x3 ../JNW_TR_SKY130A
transform 1 0 3664 0 1 0
box 3664 0 8136 3440
use JNWTR_RPPO16 x4 ../JNW_TR_SKY130A
transform 1 0 0 0 1 4040
box 0 4040 4472 7480
use JNWTR_RPPO16 x5 ../JNW_TR_SKY130A
transform 1 0 5152 0 1 4040
box 5152 4040 9624 7480
use JNWATR_PCH_4C5F0 x5[3:0] ../JNW_ATR_SKY130A
transform 1 0 10304 0 1 4040
box 10304 4040 11456 4840
use JNWATR_PCH_4C5F0 x5[3:0] ../JNW_ATR_SKY130A
transform 1 0 10304 0 1 4840
box 10304 4840 11456 5640
use JNWATR_PCH_4C5F0 x5[3:0] ../JNW_ATR_SKY130A
transform 1 0 10304 0 1 5640
box 10304 5640 11456 6440
use JNWATR_PCH_4C5F0 x5[3:0] ../JNW_ATR_SKY130A
transform 1 0 10304 0 1 6440
box 10304 6440 11456 7240
use JNWATR_NCH_4C5F0 x6 ../JNW_ATR_SKY130A
transform 1 0 12136 0 1 4040
box 12136 4040 13288 4840
use JNWATR_PCH_4C5F0 x6[3:0] ../JNW_ATR_SKY130A
transform 1 0 13968 0 1 4040
box 13968 4040 15120 4840
use JNWATR_PCH_4C5F0 x6[3:0] ../JNW_ATR_SKY130A
transform 1 0 13968 0 1 4840
box 13968 4840 15120 5640
use JNWATR_PCH_4C5F0 x6[3:0] ../JNW_ATR_SKY130A
transform 1 0 13968 0 1 5640
box 13968 5640 15120 6440
use JNWATR_PCH_4C5F0 x6[3:0] ../JNW_ATR_SKY130A
transform 1 0 13968 0 1 6440
box 13968 6440 15120 7240
use JNWATR_NCH_4C5F0 x7 ../JNW_ATR_SKY130A
transform 1 0 15800 0 1 4040
box 15800 4040 16952 4840
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 16952 7480
<< end >>
