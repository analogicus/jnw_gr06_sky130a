magic
tech sky130A
magscale 1 2
timestamp 1742943600
<< checkpaint >>
rect 0 0 2304 800
use JNWATR_PCH_4C5F0 x1 ../JNW_ATR_SKY130A
transform 1 0 0 0 1 0
box 0 0 1152 800
use JNWATR_PCH_4C5F0 x2 ../JNW_ATR_SKY130A
transform 1 0 1152 0 1 0
box 1152 0 2304 800
use JNWATR_NCH_4C5F0 x3[1:0] ../JNW_ATR_SKY130A
transform 1 0 2304 0 1 0
box 2304 0 3456 800
use JNWATR_NCH_4C5F0 x3[1:0] ../JNW_ATR_SKY130A
transform 1 0 2304 0 1 800
box 2304 800 3456 1600
use JNWATR_NCH_4C5F0 x4[1:0] ../JNW_ATR_SKY130A
transform 1 0 3456 0 1 0
box 3456 0 4608 800
use JNWATR_NCH_4C5F0 x4[1:0] ../JNW_ATR_SKY130A
transform 1 0 3456 0 1 800
box 3456 800 4608 1600
use JNWATR_PCH_4C5F0 x5[3:0] ../JNW_ATR_SKY130A
transform 1 0 4608 0 1 0
box 4608 0 5760 800
use JNWATR_PCH_4C5F0 x5[3:0] ../JNW_ATR_SKY130A
transform 1 0 4608 0 1 800
box 4608 800 5760 1600
use JNWATR_PCH_4C5F0 x5[3:0] ../JNW_ATR_SKY130A
transform 1 0 4608 0 1 1600
box 4608 1600 5760 2400
use JNWATR_PCH_4C5F0 x5[3:0] ../JNW_ATR_SKY130A
transform 1 0 4608 0 1 2400
box 4608 2400 5760 3200
use JNWATR_PCH_4C5F0 x6[3:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 0
box 5760 0 6912 800
use JNWATR_PCH_4C5F0 x6[3:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 800
box 5760 800 6912 1600
use JNWATR_PCH_4C5F0 x6[3:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 1600
box 5760 1600 6912 2400
use JNWATR_PCH_4C5F0 x6[3:0] ../JNW_ATR_SKY130A
transform 1 0 5760 0 1 2400
box 5760 2400 6912 3200
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 2304 800
<< end >>
