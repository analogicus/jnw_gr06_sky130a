magic
tech sky130A
timestamp 1742998585
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 7284 0 1 2400
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1734044400
transform 1 0 7284 0 1 2000
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1734044400
transform 1 0 7284 0 1 1600
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1734044400
transform 1 0 7284 0 1 800
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1734044400
transform 1 0 7284 0 1 400
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1734044400
transform 1 0 7284 0 1 0
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2
timestamp 1734044400
transform 1 0 3916 0 1 0
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa3
timestamp 1734044400
transform 1 0 3920 0 1 400
box -92 -64 668 464
use JNWTR_RPPO16  xb5 ../JNW_TR_SKY130A
timestamp 1742987017
transform 1 0 4752 0 1 1759
box 0 0 2236 1720
use JNWTR_RPPO16  xc4
timestamp 1742987017
transform 1 0 4756 0 1 0
box 0 0 2236 1720
use JNWTR_RPPO16  xd3
timestamp 1742987017
transform 1 0 4760 0 1 -1832
box 0 0 2236 1720
use JNWATR_PCH_4C5F0  xe5[3:0]
timestamp 1734044400
transform 1 0 7284 0 1 1200
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xe6[3:0]
timestamp 1734044400
transform 1 0 7284 0 1 2800
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xf6 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 8134 0 1 0
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xf7
timestamp 1734044400
transform 1 0 8130 0 1 400
box -92 -64 668 464
<< properties >>
string FIXED_BBOX 0 0 8436 1720
<< end >>
