magic
tech sky130A
magscale 1 2
timestamp 1743272310
<< locali >>
rect 13014 17362 13254 19656
rect 13014 17122 20142 17362
rect 11348 16956 11724 17068
rect 13014 16804 13254 17122
rect 10082 16564 10222 16804
rect 12880 16564 13254 16804
rect 16708 14412 16900 14640
rect 17732 14412 17924 14640
rect 16708 14404 17942 14412
rect 16708 14248 17098 14404
rect 17254 14248 17942 14404
rect 16708 14220 17942 14248
rect 17742 13546 17934 14220
rect 13852 13354 17934 13546
rect 10020 12426 10160 12666
rect 10794 12426 10920 12666
rect 11148 12426 11160 12666
rect 11436 9616 11676 9622
rect 11436 9388 11442 9616
rect 11670 9388 11676 9616
rect 11436 9344 11676 9388
rect 11288 9104 11676 9344
rect 11436 8456 11676 9104
rect 11306 5757 11676 8456
rect 13852 2914 14044 13354
rect 17742 13314 17934 13354
rect 19902 13250 20142 17122
rect 18690 2914 22122 4842
rect 12058 1706 22122 2914
rect 12058 1644 19410 1706
<< viali >>
rect 13014 19656 13254 19884
rect 9854 16564 10082 16804
rect 10942 16570 11170 16798
rect 11968 16564 12196 16804
rect 17098 14248 17254 14404
rect 9792 12426 10020 12666
rect 10920 12426 11148 12666
rect 11442 9388 11670 9616
<< metal1 >>
rect 10292 19884 13266 19890
rect 10292 19656 13014 19884
rect 13254 19656 13266 19884
rect 10292 19650 13266 19656
rect 14726 17698 14918 17704
rect 10104 17506 14726 17698
rect 14726 17500 14918 17506
rect 9848 16804 10088 16816
rect 11962 16804 12202 16816
rect 9054 16564 9854 16804
rect 10082 16564 10088 16804
rect 10930 16798 11968 16804
rect 10930 16570 10942 16798
rect 11170 16570 11968 16798
rect 10930 16564 11968 16570
rect 12196 16564 12202 16804
rect 9054 13328 9294 16564
rect 9848 16552 10088 16564
rect 11962 16552 12202 16564
rect 16964 15180 17028 16706
rect 17348 15248 17540 15254
rect 17348 15050 17540 15056
rect 17092 14404 17260 14696
rect 17092 14248 17098 14404
rect 17254 14248 17260 14404
rect 17092 14236 17260 14248
rect 12362 13328 12602 13334
rect 9054 13088 12362 13328
rect 9054 12666 9294 13088
rect 12362 13082 12602 13088
rect 9786 12666 10026 12678
rect 9054 12426 9792 12666
rect 10020 12426 10026 12666
rect 9054 12410 9294 12426
rect 9786 12414 10026 12426
rect 10914 12666 11154 12678
rect 10914 12426 10920 12666
rect 11148 12426 11676 12666
rect 10914 12414 11154 12426
rect 11436 9616 11676 12426
rect 11436 9388 11442 9616
rect 11670 9388 11676 9616
rect 11436 9376 11676 9388
rect 18609 8613 18675 8619
rect 18609 8384 18675 8547
rect 20591 8458 20657 8464
rect 20591 8386 20657 8392
rect 24286 6350 25414 6542
rect 2532 5414 2538 5606
rect 2730 5414 2736 5606
<< via1 >>
rect 14726 17506 14918 17698
rect 17348 15056 17540 15248
rect 12362 13088 12602 13328
rect 18609 8547 18675 8613
rect 20591 8392 20657 8458
rect 2538 5414 2730 5606
<< metal2 >>
rect 14720 17506 14726 17698
rect 14918 17506 14924 17698
rect 14726 15930 14918 17506
rect 14726 15739 14918 15748
rect 17348 15718 17540 15727
rect 17348 15248 17540 15536
rect 17342 15056 17348 15248
rect 17540 15056 17546 15248
rect 18609 13753 18675 13762
rect 12411 13328 17427 13343
rect 12356 13088 12362 13328
rect 12602 13140 17427 13328
rect 12602 13088 12608 13140
rect 13889 11697 14092 13140
rect 13889 11494 18356 11697
rect 18153 8370 18356 11494
rect 18609 8613 18675 13697
rect 18603 8547 18609 8613
rect 18675 8547 18681 8613
rect 20585 8456 20591 8458
rect 20454 8392 20591 8456
rect 20657 8392 20663 8458
rect 20454 8370 20657 8392
rect 18153 8167 20657 8370
rect 20454 8164 20656 8167
rect 2538 5606 2730 5612
rect 2538 5406 2730 5414
rect 2538 5214 2548 5406
rect 2730 5214 2739 5406
<< via2 >>
rect 14726 15748 14918 15930
rect 17348 15536 17540 15718
rect 18609 13697 18675 13753
rect 2548 5214 2730 5406
<< metal3 >>
rect 14721 15930 14923 15935
rect 14721 15748 14726 15930
rect 14918 15748 14923 15930
rect 14721 15743 14923 15748
rect 14726 14896 14918 15743
rect 15990 15531 15996 15723
rect 16186 15718 17545 15723
rect 16186 15536 17348 15718
rect 17540 15536 17545 15718
rect 16186 15531 17545 15536
rect 15297 13758 15363 14397
rect 15297 13753 18680 13758
rect 15297 13697 18609 13753
rect 18675 13697 18680 13753
rect 15297 13692 18680 13697
rect 2543 5406 2735 5411
rect 2543 5214 2548 5406
rect 2730 5214 2966 5406
rect 3156 5214 3162 5406
rect 2543 5209 2735 5214
<< via3 >>
rect 15996 15531 16186 15723
rect 2966 5214 3156 5406
<< metal4 >>
rect 15995 15723 16187 15724
rect 15400 15531 15996 15723
rect 16186 15531 16187 15723
rect 15400 14904 15592 15531
rect 15995 15530 16187 15531
rect 3696 5544 4346 5736
rect 2965 5406 3157 5407
rect 3696 5406 3888 5544
rect 2965 5214 2966 5406
rect 3156 5214 3888 5406
rect 2965 5213 3157 5214
use JNWATR_PCH_2C1F2  JNWATR_PCH_2C1F2_0 JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 16804 0 1 14488
box -184 -128 1208 928
use JNWTR_CAPX1  JNWTR_CAPX1_1 JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 14660 0 1 14036
box 0 0 1080 1080
use JNWTR_RPPO4  JNWTR_RPPO4_0 JNW_TR_SKY130A
timestamp 1743265964
transform 1 0 9596 0 1 13644
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_1
timestamp 1743265964
transform 1 0 11604 0 1 13644
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_2
timestamp 1743265964
transform 1 0 9532 0 1 9506
box 0 0 1880 3440
use OTA  OTA_0
timestamp 1743272310
transform 1 0 13972 0 1 2970
box 0 -480 10506 10458
use temp_affected_current  temp_affected_current_0
timestamp 1743272310
transform 1 0 3384 0 1 6522
box -9440 -4968 8788 13334
<< labels >>
flabel space 21642 6350 24958 6542 0 FreeSans 1600 0 0 0 OUT
port 1 nsew
flabel space 3265 12106 3692 19835 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel space -1092 1652 7684 3310 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal1 16964 16642 17028 16706 0 FreeSans 1600 0 0 0 reset
port 5 nsew
flabel space 6686 1658 12118 3424 0 FreeSans 1600 0 0 0 VSS
port 6 nsew
flabel metal1 25222 6350 25414 6542 0 FreeSans 1600 0 0 0 OUT
port 7 nsew
flabel space 3242 19638 4830 19830 0 FreeSans 1600 0 0 0 VDD
port 8 nsew
<< end >>
