magic
tech sky130A
magscale 1 2
timestamp 1743679690
<< locali >>
rect 17256 11684 33115 13304
rect 21942 11590 33115 11684
rect 26800 11104 27012 11110
rect 26800 10904 26806 11104
rect 27006 10904 27012 11104
rect -788 526 178 10894
rect 26800 10694 27012 10904
rect 26794 10462 27012 10694
rect 10902 6316 15356 6732
rect 11558 1638 12366 2946
rect 13286 2788 17710 3118
rect 17446 1638 17730 2788
rect 11558 1420 17730 1638
rect -788 364 5020 526
rect 11558 382 12366 1420
rect 17446 382 17730 1420
rect -788 266 8426 364
rect 11558 266 17730 382
rect -788 -82 17826 266
rect 20212 -82 20610 10144
rect 26794 10014 27006 10462
rect 25470 -82 28700 1514
rect -788 -527 29754 -82
rect 31401 -527 33115 11590
rect -788 -2241 33115 -527
rect -788 -2274 29754 -2241
rect -782 -2330 29754 -2274
rect -782 -2344 24 -2330
<< viali >>
rect 26806 10904 27006 11104
<< metal1 >>
rect -758 16836 30020 19068
rect -746 11268 9880 16836
rect 7032 10754 9872 11268
rect 8406 9136 9872 10754
rect 15966 9626 17074 16836
rect 21319 12621 21385 16305
rect 21313 12555 21319 12621
rect 21385 12555 21391 12621
rect 26132 11104 27028 16836
rect 26132 10904 26806 11104
rect 27006 10904 27028 11104
rect 26132 10898 27028 10904
rect 26800 10892 27012 10898
rect 15820 9464 17074 9626
rect 15820 9318 16012 9464
rect 8392 8218 11338 9136
rect 8406 5320 9872 8218
rect 19943 7465 20009 7471
rect 16581 7399 19943 7465
rect 19943 7393 20009 7399
rect 17160 6782 17604 7026
rect 25117 5457 25183 5463
rect 8406 5294 9586 5320
rect 25117 5186 25183 5391
rect 27091 5260 27157 5266
rect 27091 5188 27157 5194
rect 31908 3344 32100 3766
rect 30714 3152 32100 3344
<< via1 >>
rect 21319 12555 21385 12621
rect 19943 7399 20009 7465
rect 25117 5391 25183 5457
rect 27091 5194 27157 5260
<< metal2 >>
rect 21319 12621 21385 12627
rect 19937 7399 19943 7465
rect 20009 7399 20015 7465
rect 19943 5457 20009 7399
rect 21319 6303 21385 12555
rect 21319 6237 27157 6303
rect 19510 5391 19519 5457
rect 19575 5391 25117 5457
rect 25183 5391 25189 5457
rect 27091 5260 27157 6237
rect 27085 5194 27091 5260
rect 27157 5194 27163 5260
<< via2 >>
rect 19519 5391 19575 5457
<< metal3 >>
rect 19514 5457 19580 5462
rect 19215 5391 19519 5457
rect 19575 5391 19580 5457
rect 19215 5386 19580 5391
rect 19215 4575 19281 5386
use JNWTR_CAPX1  JNWTR_CAPX1_0 JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 18734 0 1 3742
box 0 0 1080 1080
use JNWTR_RPPO4  JNWTR_RPPO4_0 JNW_TR_SKY130A
timestamp 1743265964
transform 1 0 21466 0 1 13278
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_1
timestamp 1743265964
transform 1 0 17214 0 1 13246
box 0 0 1880 3440
use JNWTR_RPPO4  JNWTR_RPPO4_2
timestamp 1743265964
transform 1 0 19348 0 1 13262
box 0 0 1880 3440
use OTA  OTA_0
timestamp 1743679690
transform 1 0 20470 0 1 -228
box 0 -480 10506 10458
use temp_affected_current  temp_affected_current_0
timestamp 1743679690
transform 1 0 0 0 1 0
box 0 -294 23688 17114
<< labels >>
flabel locali 24 -2330 17834 -82 0 FreeSans 1600 0 0 0 VSS
port 9 nsew
flabel metal1 -758 16836 16048 19068 0 FreeSans 1600 0 0 0 VDD
port 11 nsew
flabel metal1 17160 6782 17604 7026 0 FreeSans 1600 0 0 0 reset
port 13 nsew
flabel space 28140 3152 31548 3344 0 FreeSans 1600 0 0 0 OUT
port 17 nsew
flabel metal1 31908 3152 32100 3766 0 FreeSans 1600 0 0 0 OUT
port 19 nsew
<< end >>
