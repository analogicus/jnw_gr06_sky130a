magic
tech sky130A
timestamp 1742987825
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 576 0 1 2400
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1734044400
transform 1 0 576 0 1 2000
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1734044400
transform 1 0 576 0 1 1599
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1734044400
transform 1 0 576 0 1 800
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1734044400
transform 1 0 576 0 1 400
box -92 -64 668 464
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1734044400
transform 1 0 576 0 1 0
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa2
timestamp 1734044400
transform 1 0 -381 0 1 0
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xa3
timestamp 1734044400
transform 1 0 -380 0 1 400
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xb5[3:0]
timestamp 1734044400
transform 1 0 576 0 1 1200
box -92 -64 668 464
use JNWATR_PCH_4C5F0  xb6[3:0]
timestamp 1734044400
transform 1 0 576 0 1 2800
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xc6 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 2400 0 1 -4
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xc7
timestamp 1734044400
transform 1 0 2399 0 1 400
box -92 -64 668 464
use JNWTR_RPPO16  xd5 ../JNW_TR_SKY130A
timestamp 1742987017
transform 1 0 1710 0 1 1223
box 0 0 2236 1720
use JNWTR_RPPO16  xe4
timestamp 1742987017
transform 1 0 4035 0 1 205
box 0 0 2236 1720
use JNWTR_RPPO16  xf3
timestamp 1742987017
transform 1 0 6435 0 1 688
box 0 0 2236 1720
<< properties >>
string FIXED_BBOX 0 0 8436 1720
<< end >>
